// SBOX 2 from the DES standard
module sbox2 (
    input  wire [5:0] in,   // 6-bit input
    output reg  [3:0] out   // 4-bit output
);

    wire [1:0] row;
    wire [3:0] col;

    assign row = {in[5], in[0]};
    assign col = in[4:1];

    always @(*) begin
        case ({row, col})
            6'b000000: out = 4'd15;
            6'b000001: out = 4'd1;
            6'b000010: out = 4'd8;
            6'b000011: out = 4'd14;
            6'b000100: out = 4'd6;
            6'b000101: out = 4'd11;
            6'b000110: out = 4'd3;
            6'b000111: out = 4'd4;
            6'b001000: out = 4'd9;
            6'b001001: out = 4'd7;
            6'b001010: out = 4'd2;
            6'b001011: out = 4'd13;
            6'b001100: out = 4'd12;
            6'b001101: out = 4'd0;
            6'b001110: out = 4'd5;
            6'b001111: out = 4'd10;

            6'b010000: out = 4'd3;
            6'b010001: out = 4'd13;
            6'b010010: out = 4'd4;
            6'b010011: out = 4'd7;
            6'b010100: out = 4'd15;
            6'b010101: out = 4'd2;
            6'b010110: out = 4'd8;
            6'b010111: out = 4'd14;
            6'b011000: out = 4'd12;
            6'b011001: out = 4'd0;
            6'b011010: out = 4'd1;
            6'b011011: out = 4'd10;
            6'b011100: out = 4'd6;
            6'b011101: out = 4'd9;
            6'b011110: out = 4'd11;
            6'b011111: out = 4'd5;

            6'b100000: out = 4'd0;
            6'b100001: out = 4'd14;
            6'b100010: out = 4'd7;
            6'b100011: out = 4'd11;
            6'b100100: out = 4'd10;
            6'b100101: out = 4'd4;
            6'b100110: out = 4'd13;
            6'b100111: out = 4'd1;
            6'b101000: out = 4'd5;
            6'b101001: out = 4'd8;
            6'b101010: out = 4'd12;
            6'b101011: out = 4'd6;
            6'b101100: out = 4'd9;
            6'b101101: out = 4'd3;
            6'b101110: out = 4'd2;
            6'b101111: out = 4'd15;

            6'b110000: out = 4'd13;
            6'b110001: out = 4'd8;
            6'b110010: out = 4'd10;
            6'b110011: out = 4'd1;
            6'b110100: out = 4'd3;
            6'b110101: out = 4'd15;
            6'b110110: out = 4'd4;
            6'b110111: out = 4'd2;
            6'b111000: out = 4'd11;
            6'b111001: out = 4'd6;
            6'b111010: out = 4'd7;
            6'b111011: out = 4'd12;
            6'b111100: out = 4'd0;
            6'b111101: out = 4'd5;
            6'b111110: out = 4'd14;
            6'b111111: out = 4'd9;

            default: out = 4'd0;
        endcase
    end

endmodule
